module main

import time

fn main() {
	mut game := new_game()
	game.g.run()
}

// Disables vsync, but only works on linux
@[if linux]
fn C._sapp_glx_swapinterval(int)

// frame gets called everytime a new frame is drawn to the screen.
fn frame(mut game Game) {
	game.current_time = time.now().unix_milli()
	game.delta_time = game.current_time - game.last_time
	game.last_time = game.current_time

	game.update()
	game.g.begin()
	game.draw()
	game.g.end()
}
